`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:58:01 06/03/2017 
// Design Name: 
// Module Name:    Memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Memory(
    input MemRead,
    input MemWrite,
    input [31:0] Address,
    input [31:0] WriteData,
	 input newchar,
	 input [15:0] char,
    output reg [31:0] MemData,
	 output wire [31:0] a3
    );

	reg [31:0] block [0:499];
	assign a3 = block[7];
	
	reg [1:0] contador = 0; //se utiliza para saber si viene operacion, num1 o num2

	integer i = 0;
	initial begin 
		for (i=91;i<500;i=i+1) begin
			block[i] <= 32'b0;
		end
		MemData <= 32'b0;
		block[38] <= 32'b00100000000010110000000000000001;
		block[39] <= 32'b00100000000011000000000000000010;
		block[40] <= 32'b00100000000011010000000000000011;
		block[41] <= 32'b00100000000011100000000000000100;
		block[42] <= 32'b00100000000011110000000000000101;
		block[43] <= 32'b00100000000100000000000000000110;
		block[44] <= 32'b00100000000100010000000000000111;
		block[45] <= 32'b00100000000100100000000000001000;
		block[46] <= 32'b00100000000100110000000000001001;
		block[47] <= 32'b00100000000101000000000000001010;
		block[49] <= 32'b00100000000101010000000000001011;
		block[50] <= 32'b00100000000101100000000000001100;
		block[51] <= 32'b00100000000101110000000000001101;
		block[52] <= 32'b10001100000001100000000000100011;
		block[53] <= 32'b00010000000001101111111111111110;
		block[54] <= 32'b00110000000001110000000000000000;
		block[55] <= 32'b10001100000010000000000000100100;
		block[56] <= 32'b00010001000000001111111111111110;
		block[57] <= 32'b10001100000001000000000000100001;
		block[58] <= 32'b10001100000010010000000000100101;
		block[59] <= 32'b00010001001000001111111111111110;
		block[60] <= 32'b10001100000001010000000000100010;
		block[61] <= 32'b10101100000000000000000000100100;
		block[62] <= 32'b00010001011001100000000000001111;
		block[63] <= 32'b00010001100001100000000000010000;
		block[64] <= 32'b00010001101001100000000000010011;
		block[65] <= 32'b00010001110001100000000000100001;
		block[66] <= 32'b00010001111001100000000000101001;
		block[67] <= 32'b00010010000001100000000000101000;
		block[68] <= 32'b00010010001001100000000000100111;
		block[69] <= 32'b00010010010001100000000000101000;
		block[70] <= 32'b00010010011001100000000000101001;
		block[71] <= 32'b00010010100001100000000000101010;
		block[72] <= 32'b00010010101001100000000000101100;
		block[73] <= 32'b00010010110001100000000000101101;
		block[74] <= 32'b00010010111001100000000000101100;
		block[75] <= 32'b10101100000000000000000000100011;
		block[76] <= 32'b10101100000000000000000000100101;
		block[77] <= 32'b00001000000000000000000000001101;
		block[78] <= 32'b00000000100001010011100000100000;
		block[79] <= 32'b00001000000000000000000001010111;
		block[80] <= 32'b00000000101000000010100000100111;
		block[81] <= 32'b00100000101001010000000000000001;
		block[82] <= 32'b00000000100001010011100000100000;
		block[83] <= 32'b00001000000000000000000001010111;
		block[84] <= 32'b00100000000000100000000000000000;
		block[85] <= 32'b00100000000010000000000000000001;
		block[86] <= 32'b00100000000010010000000000000000;
		block[87] <= 32'b00010000101000000000000000001001;
		block[88] <= 32'b00000001000001010100100000100100;
		block[89] <= 32'b00100000000000010000000000000001;
		block[90] <= 32'b00010000001010010000000000000010;
		block[91] <= 32'b00100000000000010000000000000000;
		block[92] <= 32'b00010000001010010000000000000001;
		block[93] <= 32'b00000000010001000001000000100000;
		block[94] <= 32'b00000000000001000010000001000000;
		block[95] <= 32'b00000000000001010010100001000010;
		block[96] <= 32'b00001000000000000000000000110000;
		block[97] <= 32'b00100000010001110000000000000000;
		block[98] <= 32'b00001000000000000000000001010111;
		block[99] <= 32'b00000000000001000100000000100000;
		block[100] <= 32'b00100000000010100000000000000000;
		block[101] <= 32'b00000001000001010100000000100010;
		block[102] <= 32'b00100001010010100000000000000001;
		block[103] <= 32'b00000001000001010101100000101010;
		block[104] <= 32'b00010101011000000000000000000001;
		block[105] <= 32'b00001000000000000000000000111110;
		block[106] <= 32'b00100001010001110000000000000000;
		block[107] <= 32'b00001000000000000000000001010111;
		block[108] <= 32'b00000000100001010011100000100100;
		block[109] <= 32'b00001000000000000000000001010111;
		block[110] <= 32'b00000000100001010011100000100101;
		block[111] <= 32'b00001000000000000000000001010111;
		block[112] <= 32'b00000000100000000011100000100111;
		block[113] <= 32'b00001000000000000000000001010111;
		block[114] <= 32'b00000000100001010011100000100100;
		block[115] <= 32'b00000000111000000011100000100111;
		block[116] <= 32'b00001000000000000000000001010111;
		block[117] <= 32'b00000000100001010011100000100111;
		block[118] <= 32'b00001000000000000000000001010111;
		block[119] <= 32'b00000000100001010100000000100100;
		block[120] <= 32'b00000001000000000100000000100111;
		block[121] <= 32'b00000000100001010011100000100101;
		block[122] <= 32'b00000000111010000011100000100100;
		block[123] <= 32'b00010010111001100000000000000001;
		block[124] <= 32'b00001000000000000000000001010111;
		block[125] <= 32'b00000000111000000011100000100111;
		block[126] <= 32'b10101100000000000000000000100011;
		block[127] <= 32'b10101100000000000000000000100101;
		block[128] <= 32'b00100000000010100000000000000001;
		block[129] <= 32'b00001000000000000000000000001101;
		
	end

	always @ (*) begin
		if (newchar)
			if (char[15:8] != 8'hF0) begin
				contador = contador + 1;
				if (contador == 0) begin
					block[35] <= {24'b000000000000000000000000,char[7:0]};
				end
				else if (contador == 1) begin
					block[33] <= {24'b000000000000000000000000,char[7:0]};
					block[36] <= 1;
				end
				else if (contador == 2) begin
					block[34] <= {24'b000000000000000000000000,char[7:0]};
					block[37] <= 1;
				end
			end
		else
			begin
				if (MemRead)
					MemData <= block[Address];
				else if (MemWrite)
					block[Address] <= WriteData;
				else
					MemData <= 32'b0;
			end
	end

endmodule
