`timescale 1ns / 1ps
module InstructionMemory(
    output reg[31:0] RA, /* Read Data Output*/
    input [31:0] A /* Adress */
    );

	always @ (*) begin
		case (A)
			32'h00000004: RA = 32'hE3A00000; //MOV		R0, #0x0
			32'h00000008: RA = 32'hE3A04004; //MOV		R4, #0x00000004
			32'h0000000c: RA = 32'hE3A05010; //MOV		R5, #0x00000010
			32'h00000010: RA = 32'hE3A06014; //MOV		R6, #0x00000014
			32'h00000014: RA = 32'hE3A07018; //MOV		R7, #0x00000018
			23'h00000018: RA = 32'hE3A0D024; //MOV		R13, OPA
			32'h0000001c: RA = 32'hE3A0801C; //MOV		R8, #0x0000001c
			//HEPHAESTUS
			32'h00000020: RA = 32'hEAFFFFFE; //B		HEPHAESTUS
			//OPA
			32'h00000024: RA = 32'hE5941000; //LDR		R1, [R4, R0] 
			32'h00000028: RA = 32'hE351000A; //CMP		R1, #10
			32'h0000002c: RA = 32'hAA000006; //BGE		SAVEOP
			32'h00000030: RA = 32'hE5952000; //LDR		R2, [R5, #0] 
			32'h00000034: RA = 32'hE1A03182; //LSL		R3, R2, #3
			32'h00000038: RA = 32'hE1A02082; //LSL		R2, R2, #1
			32'h0000003c: RA = 32'hE0822003; //ADD		R2, R2, R3
			32'h00000040: RA = 32'hE0822001; //ADD		R2, R2, R1
			32'h00000044: RA = 32'hE5852000; //STR		R2, [R5, #0]
			32'h00000048: RA = 32'hEAFFFFF4; //B		HEPHAESTUS
			//SAVEOP
			32'h0000004c: RA = 32'hE7871000; //STR		R1, [R7, R0]
			32'h00000050: RA = 32'hE3A0D058; //MOV		R13, #17
			32'h00000054: RA = 32'hEAFFFFF1; //B		HEPHAESTUS
			//OPB
			32'h00000058: RA = 32'hE7941000; //LDR		R1, [R4, R0]
			32'h0000005c: RA = 32'hE351000F; //CMP		R1, #15
			32'h00000060: RA = 32'h0A000006; //BEQ		EXE
			32'h00000064: RA = 32'hE7962000; //LDR		R2, [R6, R0]
			32'h00000068: RA = 32'hE1A03182; //LSL		R3, R2, #3
			32'h0000006c: RA = 32'hE1A02082; //LSL		R2, R2, #1
			32'h00000070: RA = 32'hE0822003; //ADD		R2, R2, R3
			32'h00000074: RA = 32'hE0822001; //ADD		R2, R2, R1
			32'h00000078: RA = 32'hE7861000; //STR		R1, [R6, R0]
			32'h0000007c: RA = 32'hEAFFFFE7; //B		HEPHAESTUS
			//EXE
			32'h00000080: RA = 32'hE7971000; //LDR		R1, [R7, R0] 
			32'h00000084: RA = 32'hE7952000; //LDR		R2, [R5, R0]
			32'h00000088: RA = 32'hE7963000; //LDR		R3, [R6, R0]
			32'h0000008c: RA = 32'hE351000A; //CMP 	R1, #10
			32'h00000090: RA = 32'h0A000007; //B 		SUM
			32'h00000094: RA = 32'hE351000B; //CMP 	R1, #11
			32'h00000098: RA = 32'h0A000007; //B		SUB
			32'h0000009c: RA = 32'hE351000C; //CMP 	R1, #12
			32'h000000a0: RA = 32'h0A000007; //B		MUL
			32'h000000a4: RA = 32'hE351000D; //CMP 	R1, #13
			32'h000000a8: RA = 32'h0A00000A; //B		DIV
			32'h000000ac: RA = 32'hE351000E; //CMP 	R1, #14
			32'h000000b0: RA = 32'h0A00000D; //B		MOD
			//SUM
			32'h000000b4: RA = 32'hE0820003; //ADD		R0, R2, R3
			32'h000000b8: RA = 32'hEA000011; //B		SAVEAN
			//SUB
			32'h000000bc: RA = 32'hE0420003; //SUB		R0, R2, R3
			32'h000000c0: RA = 32'hEA00000F; //B		SAVEAN
			//MUL
			32'h000000c4: RA = 32'hE0800002; //ADD		R0, R0, R2
			32'h000000c8: RA = 32'hE2433001; //SUB		R3, R3, #1
			32'h000000cc: RA = 32'hE3530000;	//CMP 	R3, #0
			32'h000000d0: RA = 32'h0A00000B; //BEQ		SAVEAN
			32'h000000d4: RA = 32'hEAFFFFFA; //B		MUL
			//DIV
			32'h000000d8: RA = 32'hE1520003;	//CMP 	R2, R3
			32'h000000dc: RA = 32'hBA000008;	//BLT		SAVEAN
			32'h000000e0: RA = 32'hE2800001; //ADD		R0, R0, #1
			32'h000000e4: RA = 32'hE0422003; //SUB		R2, R2, R3
			32'h000000e8: RA = 32'hEAFFFFFA; //B		DIV
			//MOD
			32'h000000ec: RA = 32'hE1520003;	//CMP 	R2, R3
			32'h000000f0: RA = 32'hB2820000;	//ADDLT	R0, R2, #0
			32'h000000f4: RA = 32'hE1520003;	//CMP 	R2, R3
			32'h000000f8: RA = 32'hBA000001;	//BLT		SAVEAN
			32'h000000fc: RA = 32'hE0422003; //SUB		R2, R2, R3
			32'h00000100: RA = 32'hEAFFFFF9; //B		MOD
			//SAVEAN
			32'h00000104: RA = 32'hE5880000; //STR		R0, [R8, #0]
			32'h00000108: RA = 32'hE3A0D120; //MOV		R13, CLEAR
			32'h0000010c: RA = 32'hEAFFFFC3; //B 		HEPHAESTUS
			//CLEAR
			32'h00000120: RA = 32'h00000000; 
			default: RA = 32'b0;
		endcase
	end

endmodule
